`timescale 1ns/1ps
// Verilog code for carry look-ahead adder
module cla_adder (in1, in2, carry_in, sum, carry_out);
parameter DATA_WID = 16;   // match testbench

input  [DATA_WID - 1:0] in1;
input  [DATA_WID - 1:0] in2;
input  carry_in;
output [DATA_WID - 1:0] sum;
output carry_out;

wire [DATA_WID - 1:0] gen;
wire [DATA_WID - 1:0] pro;
wire [DATA_WID:0] carry_tmp;

genvar j, i;
generate
    assign carry_tmp[0] = carry_in;
    
    // Carry generator
    for (j = 0; j < DATA_WID; j = j + 1) begin: carry_generator
        assign gen[j] = in1[j] & in2[j];
        assign pro[j] = in1[j] | in2[j];
        assign carry_tmp[j+1] = gen[j] | (pro[j] & carry_tmp[j]);
    end

    // Carry out
    assign carry_out = carry_tmp[DATA_WID];
    
    // Sum bits
    for (i = 0; i < DATA_WID; i = i+1) begin: sum_without_carry
        assign sum[i] = in1[i] ^ in2[i] ^ carry_tmp[i];
    end
endgenerate
endmodule
